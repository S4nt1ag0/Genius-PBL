//------------------------------------------------------------------------------
// grn
//------------------------------------------------------------------------------
// This module performs the addition of two 4-bit numbers with a carry-in and 
// produces a 4-bit sum and a carry-out.
//
// Author: Gustavo Santiago
// Date  : Maio 2025
//------------------------------------------------------------------------------

`timescale 1ns / 1ps

module grn
#(parameter DATA_WIDTH = 8)
(
    input logic clk,
    input logic seed,
    output logic [DATA_WIDTH-1:0] out
    );

    always_ff @(posedge clk) begin: get_data
        if(clk) begin
            out <= seed;
        end
    end

endmodule